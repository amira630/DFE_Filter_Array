////////////////////////////////////////////////////////////////////////////////
// Author: Amira Atef
// Design: An integrator module.
// Date: 02-11-2025
// Description: An integration stage for CIC filter
////////////////////////////////////////////////////////////////////////////////

module INTEG #(
    parameter int DATA_WIDTH = 32'd16   , 
    parameter int ACC_WIDTH = 32'd20
) (
    input  logic                                clk         ,
    input  logic                                rst_n       ,   
    input  logic                                valid_in    ,
    input  logic signed [DATA_WIDTH - 1 : 0]    intg_in     ,
    output logic signed [ACC_WIDTH - 1 : 0]     intg_out
);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            intg_out <= {ACC_WIDTH{1'sb0}};
        end else if (valid_in) begin
            intg_out <= $signed({{(ACC_WIDTH - DATA_WIDTH){intg_in[DATA_WIDTH - 1]}}, intg_in}) + intg_out;
        end
    end
endmodule