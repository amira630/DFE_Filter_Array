module top_tb ();

    // DUT Parameters
    parameter DATA_WIDTH = 16;
    parameter DATA_FRAC  = 15;
    parameter Q = 1;
    parameter N = 1;

    // Testbench Parameters
    localparam MAX_DEC_FACTOR = 16;
    localparam DEC_WIDTH = $clog2(MAX_DEC_FACTOR);

    parameter N_SAMPLES_I   = 32000                     ;
    parameter FREQ_CLK      = 9_000_000                ;
    parameter T_CLK         = 1_000_000_000 / FREQ_CLK  ;
    parameter TOLERANCE     = 1                         ;  // Tolerance for comparison (in LSBs)

    // Signals for monitoring output
    integer                     i                                           ;
    integer                     j                                           ;
    integer                     number_of_output_samples                    ;
    integer                     total_tests                                 ;
    integer                     passed_tests                                ;
    
    real                        input_sig                                   ;
    real                        output_sig                                  ;
    real                        output_sig_exp                              ;
    
    logic [DATA_WIDTH - 1 : 0]  input_samples        [N_SAMPLES_I - 1 : 0]  ;
    logic [DATA_WIDTH - 1 : 0]  output_exp_samples   [(N_SAMPLES_I) - 1 : 0]  ;

    // DUT Signals
    logic                           clk         ;
    logic                           rst_n       ;
    logic                           valid_in    ;
    logic        [DEC_WIDTH : 0]    dec_factor  ;
    logic signed [DATA_WIDTH-1:0]   cic_in      ;
    logic signed [DATA_WIDTH-1:0]   cic_out     ;
    logic                           valid_out   ;
    logic                           overflow    ;
    logic                           underflow   ;

    CIC #(
        .DATA_WIDTH(DATA_WIDTH) , 
        .DATA_FRAC(DATA_FRAC)  ,
        .Q(Q) , 
        .N(N)
    ) DUT (
        .clk        (clk)         ,
        .rst_n      (rst_n)       ,
        .valid_in   (valid_in)    ,
        .dec_factor (dec_factor)  ,  
        .cic_in     (cic_in)      ,
        .cic_out    (cic_out)     ,
        .valid_out  (valid_out)   ,   
        .overflow   (overflow)    ,
        .underflow  (underflow) 

    );

    initial begin
        clk = 0;
        forever #(T_CLK/2) clk = ~clk;
    end

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            output_sig <= 0;
        end else if (valid_out) begin
            output_sig <= $itor($signed(cic_out)) / 32768.0;
        end
    end

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            output_sig_exp <= 0;
            j <= 0;
        end else if (valid_out) begin
            output_sig_exp <= $itor($signed(output_exp_samples[j])) / 32768.0;
            j <= j + 1;
        end
    end

    // Self-checking logic with display messages
    always @(posedge clk) begin
        if (valid_in) begin
            if ((output_sig == output_sig_exp)) begin
                passed_tests = passed_tests + 1;
                total_tests = total_tests + 1;
            end else begin
                total_tests = total_tests + 1;
                $display("[%0t]: Mismatch: Expected = %f, Got = %f", $time, output_sig_exp, output_sig);
            end
        end
    end

    initial begin
        $display("================================================================================");
        $display("                     CIC Filter Testbench Started");
        $display("================================================================================");
        $display("Configuration:");
        $display("  DATA_WIDTH = %0d, DATA_FRAC = %0d, Q = %0d, N = %0d", DATA_WIDTH, DATA_FRAC, Q, N);
        $display("  N_SAMPLES = %0d, CLK_FREQ = %0d Hz", N_SAMPLES_I, FREQ_CLK);
        $display("  TOLERANCE = %0d LSBs", TOLERANCE);
        $display("================================================================================\n");

        total_tests = 0;
        passed_tests = 0;

        // Test 1: Decimation Factor = 1 (checking disabled)
        dec_factor = 1;
        $display("\nStarting test with Decimation Factor = %0d [CHECKING DISABLED]", dec_factor);
        $display("--------------------------------------------------------------------------------");
        init();
        start_CIC();
        assert_reset();

        // Test 2: Decimation Factor = 2
        dec_factor = 8;
        $display("\nStarting test with Decimation Factor = %0d", dec_factor);
        $display("--------------------------------------------------------------------------------");
        init();
        start_CIC();
        assert_reset();

        // Test 3: Decimation Factor = 4
        dec_factor = 4;
        $display("\nStarting test with Decimation Factor = %0d", dec_factor);
        $display("--------------------------------------------------------------------------------");
        init();
        start_CIC();
        assert_reset();

        // Test 4: Decimation Factor = 8
        dec_factor = 8;
        $display("\nStarting test with Decimation Factor = %0d", dec_factor);
        $display("--------------------------------------------------------------------------------");
        init();
        start_CIC();
        assert_reset();

        // Test 5: Decimation Factor = 16
        dec_factor = 16;
        $display("\nStarting test with Decimation Factor = %0d", dec_factor);
        $display("--------------------------------------------------------------------------------");
        init();
        start_CIC();
       
        repeat (5) @(negedge clk);

        // Final summary
        $display("\n================================================================================");
        $display("                          Test Summary");
        $display("================================================================================");
        $display("Total Tests Run    : %0d", total_tests);
        $display("Tests Passed       : %0d", passed_tests);
        $display("Tests Failed       : %0d", total_tests - passed_tests);
        $display("Pass Rate          : %.2f%%", (passed_tests * 100.0) / total_tests);
        $display("================================================================================");
        
        if (passed_tests == total_tests) begin
            $display("\n*** ALL TESTS PASSED ***\n");
        end else begin
            $display("\n*** SOME TESTS FAILED ***\n");
        end

        $stop;
    end

    task init ();
        $display("  Loading input samples from input_wave.txt...");
        $readmemb("input_wave.txt", input_samples);
        assert_reset();

        if(dec_factor == 1) begin
            $display("  Loading expected output from output_D1_wave_exp.txt...");
            $readmemb("output_D1_wave_exp.txt", output_exp_samples);
        end else if (dec_factor == 2) begin
            $display("  Loading expected output from output_D2_wave_exp.txt...");
            $readmemb("output_D2_wave_exp.txt", output_exp_samples);
        end else if (dec_factor == 4) begin
            $display("  Loading expected output from output_D4_wave_exp.txt...");
            $readmemb("output_D4_wave_exp.txt", output_exp_samples);
        end else if (dec_factor == 8) begin
            $display("  Loading expected output from output_D8_wave_exp.txt...");
            $readmemb("output_D8_wave_exp.txt", output_exp_samples);
        end else if (dec_factor == 16) begin
            $display("  Loading expected output from output_D16_wave_exp.txt...");
            $readmemb("output_D16_wave_exp.txt", output_exp_samples);
        end else begin
            $display("  Loading expected output from output_wave_exp.txt...");
            $readmemb("output_wave_exp.txt", output_exp_samples);
        end
        
        rst_n      = 1;
        cic_in     = 'd0;
        valid_in   = 1'b0;
        
        repeat (1) @(negedge clk);
        $display("  Initialization complete.");
    endtask

    task assert_reset ();
        $display("  Asserting reset...");
        rst_n = 0;
        repeat (5) @(negedge clk);
        rst_n = 1;
        $display("  Reset released.");
    endtask

    task start_CIC ();
        $display("  Starting CIC filter processing with %0d input samples...", N_SAMPLES_I);
        valid_in    = 1;
        rst_n       = 1;

        i = 0;

        number_of_output_samples = N_SAMPLES_I / dec_factor;

        repeat (N_SAMPLES_I ) begin
            cic_in = input_samples[i];
            input_sig = $itor($signed(input_samples[i])) / 32768.0;
            
            i = i + 1;
            @(negedge clk);
        end

        @(negedge clk);
        valid_in   = 0;
        
        // Wait for pipeline to flush
        repeat (10) @(negedge clk);
        $display("  Input processing complete. Total output samples: %0d", number_of_output_samples);
    endtask

endmodule